module frmt1(a,b,c,e);
    input a;
    input wire [7:0] b,e;
    output reg c;
endmodule