module frmt4(a, b, c);

input a; 
input b; 
output c; 
wire a;
wire b;
reg c;