module frmt1(a,b,c,e,f);
    input a;
    input wire [7:0] b,e; 
    reg e;
    output reg c;
endmodule