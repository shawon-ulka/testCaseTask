module frmt1(a,b,c);
    input a;
    input wire b;
    output reg c;
endmodule 
