module frmt5(input a, output reg f,y,
input wire b,d,
output reg c);

endmodule