module frmt3(input a,input wire b,output reg [7:0] c,d);

endmodule