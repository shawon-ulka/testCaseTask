module frmt5(input a, output reg f,y);
input wire b,d,
inout clk;output reg name1,name2;
reg [7:0] b,d,name2,
output reg c);

endmodule