module frmt5(input a, output reg f,y);
input wire b,d,
inout clk;output reg name1,name2;
output reg c);

endmodule