module frmt2(input a,clk,be,wc
            input wire b,
            output reg c
            reg [7:0] b,
            logic c,b,a

            );
endmodule