module frmt3(input a,input wire b,output reg c);

endmodule